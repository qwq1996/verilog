`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/04/02 15:20:44
// Design Name: 
// Module Name: Temperature_controller
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Temperature_controller(
    input CLK,              //20MHz
    input rst_n,
    input Cooling,
    input [15:0] Targer_Temp,
    input CMOS_Temp_en,
    input [15:0] CMOS_Temp,
    output read_cmos_temp,
    output reg [7:0] Cooling_state ,
    output [11:0] v_monitor,
    output DAC_CS,
    output DAC_SCK,
    output DAC_SDI,
    input CLK_RST_N,
    input [63:0] SN_number,
    
    input [23:0] PID_Parameter
    );
 
/***********************************************************************************************************/
/*************************************  Start Parameter Declaration  ***************************************/
/***********************************************************************************************************/
   
/***********************************************************************************************************/
/***************************************  End Parameter Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/******************************************  Start Wire Declaration  ***************************************/
/***********************************************************************************************************/

    wire [3:0] du_reg;
    
/*************************************************************************************************************/
/*****************************************  End Wire Declaration  ********************************************/
/*************************************************************************************************************/

/***********************************************************************************************************/
/*************************************  Start Registers Declaration  ***************************************/
/***********************************************************************************************************/
    reg Cooling_state = 8'h0;
/***********************************************************************************************************/
/***************************************  End Registers Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/*****************************************  Start instants Declaration  ************************************/
/***********************************************************************************************************/
    PID_controller PID_controller_inst(
    .CLK(CLK),              //20MHz
    .rst_n(rst_n),
    .CLK_RST_N(CLK_RST_N),
    .Targer_Temp(Targer_Temp),
    .CMOS_Temp_en(CMOS_Temp_en),
    .CMOS_Temp(CMOS_Temp),
    .read_cmos_temp(read_cmos_temp),
    .du_reg(du_reg),
    .PID_Parameter(PID_Parameter)
    );
    
    TEC_controller TEC_controller_inst(
    .CLK(CLK),
    .rst_n(rst_n),
    .du_reg(du_reg),
    .Cooling(Cooling),
    .DAC_CS(DAC_CS),
    .DAC_SCK(DAC_SCK),
    .DAC_SDI(DAC_SDI),
    .v_monitor(v_monitor)
    );
/***********************************************************************************************************/
/****************************************  End of instants Declaration  ************************************/
/***********************************************************************************************************/

/*************************************************************************************************************/
/*********************************  Start Design RTL Description  ********************************************/
/*************************************************************************************************************/
        
    always@(posedge CLK)
    begin
        if(Cooling == 8'h0) Cooling_state <= 8'h0;
        else if(CMOS_Temp_en) begin
            if((Targer_Temp == CMOS_Temp) || (Targer_Temp == (CMOS_Temp + 1'b1)) || (Targer_Temp == (CMOS_Temp - 1'b1))) Cooling_state <= 8'h2;
            else Cooling_state <= 8'h1;
        end
    end
    


/*************************************************************************************************************/
/***********************************  End Design RTL Description  ********************************************/
/*************************************************************************************************************/

/*************************************************************************************************************/
/***********************************  Start test Description  ************************************************/
/*************************************************************************************************************/

//    ila_6 ila_6(
//    .clk(CLK),
//    .probe0(Targer_Temp),
//    .probe1(CMOS_Temp),
//    .probe2(Targer_Temp),
//    .probe3(SN_number)
//    );

/*************************************************************************************************************/
/*************************************  end test Description  ************************************************/
/*************************************************************************************************************/

endmodule
