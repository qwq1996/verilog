///////////////////////////////////////////////
//author:qh
//data	:20210318;
//aim	 control pwm and power to fan.
///////////////////////////////////////////////

//00->second-line   01->three-line   10->four-line
module fan_4line(
    input clk,
    input [1:0] pwm_choice,
    input [1:0] power_choice,
    input [1:0] line_choice,
    input fan_switch,
    input [11:0] freq,
    output wire pwm_out,
    output wire power_out
);
/***********************************************************************************************************/
/*************************************  Start Parameter Declaration  ***************************************/
/***********************************************************************************************************/
parameter speed_25=2'b00,speed_25_cnt=12'h080;
parameter speed_50=2'b01,speed_50_cnt=12'h100;
parameter speed_75=2'b10,speed_75_cnt=12'h200;
parameter speed_100=2'b11,speed_100_cnt=12'h400;
/***********************************************************************************************************/
/***************************************  End Parameter Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/******************************************  Start Wire Declaration  ***************************************/
/***********************************************************************************************************/

/*************************************************************************************************************/
/*****************************************  End Wire Declaration  ********************************************/
/*************************************************************************************************************/

/***********************************************************************************************************/
/*************************************  Start Registers Declaration  ***************************************/
/***********************************************************************************************************/
reg pwm;
reg power;

reg [11:0] freq_cnt=12'b0;

reg [1:0] pwm_SM=2'b0;
reg [1:0] power_SM=2'b0;

reg [11:0] mode_cnt=12'b0;

reg mode_pwm_25=1'b0;
reg mode_power_25=1'b0;

reg mode_pwm_50=1'b0;
reg mode_power_50=1'b0;

reg mode_pwm_75=1'b0;
reg mode_power_75=1'b0;
/***********************************************************************************************************/
/***************************************  End Registers Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/*****************************************  Start instants Declaration  ************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/****************************************  End of instants Declaration  ************************************/
/***********************************************************************************************************/

/*************************************************************************************************************/
/*********************************  Start Design RTL Description  ********************************************/
/*************************************************************************************************************/
assign pwm_out = fan_switch ? pwm : 1'b0;
assign power_out = fan_switch ? power : 1'b0;

always @(posedge clk)
begin
    if(mode_cnt==speed_100_cnt)
        begin
            mode_cnt<=12'b0;
        end
    else
        begin
            mode_cnt<=mode_cnt+1;
        end
end

always @(posedge clk)
begin
    power_SM<=power_choice;

    case (power_SM)
        speed_100:begin
        power<=1'b1;
        end

        speed_75:begin
        power<=mode_power_75;
        end

        speed_50:begin
        power<=mode_power_50;
        end

        speed_25:begin
        power<=mode_power_25;
        end

        default:begin
            power_SM <= speed_50;
        end
    endcase
end

always @(posedge clk)
begin
    if(line_choice==2'b00)
        begin
            pwm=1'b0;
        end
    else
        begin
        pwm_SM<=pwm_choice;
  
        case (pwm_SM)
            speed_100:begin
            pwm<=1'b1;
            end

            speed_75:begin
            pwm<=mode_pwm_75;
            end

            speed_50:begin
            pwm<=mode_pwm_50;
            end

            speed_25:begin
            pwm<=mode_pwm_25;
            end

            default:begin
                pwm_SM <= mode_pwm_50;
            end
            endcase
        end
end 

always @(posedge clk)
begin
    if(mode_cnt<=speed_75_cnt)
        begin
            mode_power_75<=1'b1;
            mode_pwm_75<=1'b1;
        end
    else
        begin
            mode_power_75<=1'b0;
            mode_pwm_75<=1'b0;
        end
end
                       
always @(posedge clk)
begin
    if(mode_cnt<=speed_50_cnt)
        begin
            mode_power_50<=1'b1;
            mode_pwm_50<=1'b1;
        end
    else
        begin
            mode_power_50<=1'b0;
            mode_pwm_50<=1'b0;
        end
end

always @(posedge clk)
begin
    if(mode_cnt<=speed_25_cnt)
        begin
            mode_power_25<=1'b1;
            mode_pwm_25<=1'b1;
        end
    else
        begin
            mode_power_25<=1'b0;
            mode_pwm_25<=1'b0;
        end
end

endmodule
/*************************************************************************************************************/
/***********************************  End Design RTL Description  ********************************************/
/*************************************************************************************************************/

/*************************************************************************************************************/
/***********************************  Start test Description  ************************************************/
/*************************************************************************************************************/

/*************************************************************************************************************/
/*************************************  end test Description  ************************************************/
/*************************************************************************************************************/
/////////////////////////////////////////////

