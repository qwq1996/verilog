// -----------------------------------------------------------------------------
// Author : qwq qwq1996@mail.ustc.edu.cn
// File   : 
// Create : 2021-1-22
// Editor : 
// -----------------------------------------------------------------------------


module EP6data_combo(
input  clk_100,
input  clk_20,
input  clk_200,

input  [31:0] data1,
input  data1_en,
input  [31:0] data2,
input  data2_en,
input  [31:0] data3,
input  data3_en,

output  [31:0] dataout,
output  dataout_en
);

/***********************************************************************************************************/
/*************************************  Start Parameter Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/***************************************  End Parameter Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/******************************************  Start Wire Declaration  ***************************************/
/***********************************************************************************************************/

wire data1_out_en;
wire rd_req;
wire [31:0] data1_fifo_q;
wire cmd_fb_empty;

/*************************************************************************************************************/
/*****************************************  End Wire Declaration  ********************************************/
/*************************************************************************************************************/

/***********************************************************************************************************/
/*************************************  Start Registers Declaration  ***************************************/
/***********************************************************************************************************/

reg[399:0] rd_req_reg;

/***********************************************************************************************************/
/***************************************  End Registers Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/*****************************************  Start instants Declaration  ************************************/
/***********************************************************************************************************/

cmd_fb u_cmd_fb (
  .rst(1'b0),                  // input wire rst
  .wr_clk(clk_100),            // input wire wr_clk
  .rd_clk(clk_100),            // input wire rd_clk
  .din(data1),                  // input wire [31 : 0] din
  .wr_en(data1_en),              // input wire wr_en
  .rd_en(rd_req),              // input wire rd_en
  .dout(data1_fifo_q),                // output wire [31 : 0] dout
  .full(),                // output wire full
  .empty(cmd_fb_empty),              // output wire empty
  .wr_rst_busy(),  // output wire wr_rst_busy
  .rd_rst_busy()  // output wire rd_rst_busy
);

/***********************************************************************************************************/
/****************************************  End of instants Declaration  ************************************/
/***********************************************************************************************************/

/*************************************************************************************************************/
/*********************************  Start Design RTL Description  ********************************************/
/*************************************************************************************************************/

assign dataout_en = data1_out_en || data2_en;
assign dataout = data1_out_en ? data1_fifo_q : data2_en ? data2 : 32'd0;
assign rd_req = rd_req_reg[398] && !cmd_fb_empty;
assign data1_out_en = rd_req_reg[399] && rd_req_reg [0];

always @(posedge clk_100 ) begin
	rd_req_reg[0]   <= !cmd_fb_empty;
	rd_req_reg[399:1] <= rd_req_reg[398:0];
end

/*************************************************************************************************************/
/***********************************  End Design RTL Description  ********************************************/
/*************************************************************************************************************/

// ila_0 ila_ep6 (
// 	.clk(clk_200), // input wire clk


// 	.probe0(rd_req), // input wire [0:0]  probe0  
// 	.probe1(dataout), // input wire [0:0]  probe1 
// 	.probe2(data1_out_en), // input wire [0:0]  probe2 
// 	.probe3(cmd_fb_empty), // input wire [0:0]  probe3 
// 	.probe4(dataout), // input wire [31:0]  probe4 
// 	.probe5(data1_fifo_q) // input wire [31:0]  probe5
// );

endmodule 